TOP_tb;
reg [5:0] in1_tb;
reg [5:0] in2_tb;
reg h2_tb;
reg f9_tb;
reg jk_tb;
reg j99_tb;
reg [31:0] bus_A_tb;
reg [6:0] clk_T_tb;
reg [15:0] module_Bus_B_tb;
wire wrr_898_tb;
wire jjh_tb;
wire [63:0] d877_tb;
wire [31:0] data_rd_T_tb;
wire [31:0] f459_87__tb;
wire bus__tb;

TOP UUT (
.in1 (in1_tb),
.in2 (in2_tb),
.h2 (h2_tb),
.f9 (f9_tb),
.jk (jk_tb),
.j99 (j99_tb),
.bus_A (bus_A_tb),
.clk_T (clk_T_tb),
.module_Bus_B (module_Bus_B_tb),
.wrr_898 (wrr_898_tb),
.jjh (jjh_tb),
.d877 (d877_tb),
.data_rd_T (data_rd_T_tb),
.f459_87_ (f459_87__tb),
.bus_ (bus__tb)
);
initial
begin
end


endmodule